//this is first file 
